' phase shift oscillator
.model npn npn bf=100
Vcc (vcc 0) pulse(iv=0 pv=12 rise=.01)
Rb1 (vcc b) 100k
Rb2 (b 0)   10k
Rc  (vcc c) 10k
Re  (e 0)   1k
Ce  (e 0)   5000u
Re2 (e2 0)  1k
Q1  (c b e)    npn
Q2  (vcc c e2) npn
C1  (e2 f1) .01u
C2  (f1 f2) .01u
C3  (f2 b)  .01u
Rf1 (f1 0)  10k
Rf2 (f2 0)  10k
